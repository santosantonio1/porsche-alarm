//---------------------------------
//--                             --
//--         M O D U L E         --
//--                             --
//---------------------------------

module rgb(
    output[2:0] color
);

//---------------------------------
//--                             --
//--       A S S I G N s         --
//--                             --
//---------------------------------

assign color = 3'b101;

endmodule