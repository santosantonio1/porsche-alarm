module rgb(
    output[2:0] color
);

assign color = 3'b101;

endmodule