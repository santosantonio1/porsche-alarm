module rgb(
    output[2:0] rgb
);

assign rgb = 3'b101;

endmodule